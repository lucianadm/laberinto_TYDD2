library verilog;
use verilog.vl_types.all;
entity matriz_pru is
    port(
        C0              : out    vl_logic_vector(3 downto 0);
        D_in_A          : in     vl_logic;
        D_in_B          : in     vl_logic;
        D_in_C          : in     vl_logic;
        D_in_D          : in     vl_logic;
        reset           : in     vl_logic;
        C13             : out    vl_logic;
        C12             : out    vl_logic;
        C11             : out    vl_logic;
        C10             : out    vl_logic;
        C103            : out    vl_logic;
        C102            : out    vl_logic;
        C101            : out    vl_logic;
        C100            : out    vl_logic;
        C113            : out    vl_logic;
        C112            : out    vl_logic;
        C111            : out    vl_logic;
        C110            : out    vl_logic;
        C123            : out    vl_logic;
        C122            : out    vl_logic;
        C121            : out    vl_logic;
        C120            : out    vl_logic;
        C133            : out    vl_logic;
        C132            : out    vl_logic;
        C131            : out    vl_logic;
        C130            : out    vl_logic;
        C14             : out    vl_logic_vector(3 downto 0);
        C15             : out    vl_logic_vector(3 downto 0);
        C2              : out    vl_logic_vector(3 downto 0);
        C3              : out    vl_logic_vector(3 downto 0);
        C4              : out    vl_logic_vector(3 downto 0);
        C5              : out    vl_logic_vector(3 downto 0);
        C6              : out    vl_logic_vector(3 downto 0);
        C7              : out    vl_logic_vector(3 downto 0);
        C8              : out    vl_logic_vector(3 downto 0);
        C9              : out    vl_logic_vector(3 downto 0)
    );
end matriz_pru;
